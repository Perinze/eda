module manager # (
  parameter DW = 2
)